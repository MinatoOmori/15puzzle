`define REGISTER_N 32

`define REGISTER_ADDR_W 5
`define REGISTER_DATA_W 32

`define REGISTER_WRITE_SEL_W 2
`define REGISTER_WRITE_SEL_ALU_OUT `REGISTER_WRITE_SEL_W'd0
`define REGISTER_WRITE_SEL_PC `REGISTER_WRITE_SEL_W'd1
`define REGISTER_WRITE_SEL_DMEM `REGISTER_WRITE_SEL_W'd2
