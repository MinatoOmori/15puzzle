`define DISABLE 1'b0
`define ENABLE 1'b1
