`define PC_OP_W 2

`define PC_OP_DEFAULT `PC_OP_W'd0
`define PC_OP_JAL `PC_OP_W'd1
`define PC_OP_JALR `PC_OP_W'd2
`define PC_OP_BRANCH `PC_OP_W'd3
